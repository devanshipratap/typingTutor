module fsm (
    output score_change,
    output ,
    input correct
    );

    wire sInitial, sCorrect, sWrong, sReset;

endmodule // fsm
