module scoreCounter (
    input clk,
    input reset,
    input incOrDec,
    output [3:0] score
    );

    reg 

endmodule
